module hello_world;

initial begin
    $display("Hello Verilog!");
end

endmodule
